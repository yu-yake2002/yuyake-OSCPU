//--Sun Jiru, Nanjing Uniersity--

`include "defines.v"

module excp_handler (
  
);

  
endmodule